----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:07:53 11/05/2021 
-- Design Name: 
-- Module Name:    BRAMHandler - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity BRAMHandler_CurveB_B00 is
	 Generic ( DataWidth : integer := 18);
    Port ( CLK_IN : in  STD_LOGIC;
			  ENA_IN : in STD_LOGIC;
           ADDRA_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DOA_OUT : out  STD_LOGIC_VECTOR(31 downto 0);
			  DOPA_OUT : out  STD_LOGIC_VECTOR(3 downto 0);
			  ENB_IN : in STD_LOGIC;
           ADDRB_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DIB_IN : in  STD_LOGIC_VECTOR(31 downto 0);
			  DIPB_IN : in  STD_LOGIC_VECTOR(3 downto 0));
end BRAMHandler_CurveB_B00;

architecture Behavioral of BRAMHandler_CurveB_B00 is

	signal REGCEA: STD_LOGIC := '0';
	signal RSTA: STD_LOGIC := '0';
	signal WEA : STD_LOGIC_VECTOR(3 downto 0)  := (others => '0');
	signal DIA : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DIPA : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');

	signal DOB : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DOPB : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');
	signal REGCEB: STD_LOGIC := '0';
	signal RSTB: STD_LOGIC := '0';
	signal WEB : STD_LOGIC_VECTOR(3 downto 0) := (others => '1');
	
begin

	-- RAMB16BWER: 16k-bit Data and 2k-bit Parity Configurable Synchronous Dual Port Block RAM with Optional Output Registers
   --             Spartan-6
   -- Xilinx HDL Language Template, version 14.7

   RAMB16BWER_inst00 : RAMB16BWER
   generic map (
      -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
      DATA_WIDTH_A => DataWidth,
      DATA_WIDTH_B => DataWidth,
      -- DOA_REG/DOB_REG: Optional output register (0 or 1)
      DOA_REG => 0,
      DOB_REG => 0,
      -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
      EN_RSTRAM_A => TRUE,
      EN_RSTRAM_B => TRUE,
     	-- INITP_00 to INITP_07: Initial memory contents.
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

		-- INIT_00 to INIT_3F: Initial memory contents.
		INIT_00 => X"0179015F0146012D011400FB00E200C900AF0096007D0064004B003200190000",
		INIT_01 => X"030A02F102D802BF02A6028D0274025B02420228020F01F601DD01C401AB0192",
		INIT_02 => X"049C0483046A04510438041F040503EC03D303BA03A10388036F0356033D0324",
		INIT_03 => X"062D061405FB05E205C905B00597057D0564054B05320519050004E704CE04B5",
		INIT_04 => X"07BC07A4078B0772075907400727070E06F506DC06C306AA06910678065F0646",
		INIT_05 => X"094B09320919090008E808CF08B6089D0884086B085208390820080707EE07D5",
		INIT_06 => X"0AD80ABF0AA70A8E0A750A5C0A440A2B0A1209F909E009C709AF0996097D0964",
		INIT_07 => X"0C640C4B0C320C1A0C010BE80BD00BB70B9E0B860B6D0B540B3B0B230B0A0AF1",
		INIT_08 => X"0DED0DD50DBC0DA40D8B0D730D5A0D410D290D100CF80CDF0CC60CAE0C950C7C",
		INIT_09 => X"0F750F5C0F440F2C0F130EFB0EE20ECA0EB10E990E800E680E4F0E370E1E0E06",
		INIT_0A => X"10FA10E210C910B110991081106810501038101F10070FEF0FD60FBE0FA60F8D",
		INIT_0B => X"127C1264124C1234121C120411EC11D411BB11A3118B1173115B1143112A1112",
		INIT_0C => X"13FC13E413CC13B4139C1384136C1354133C1324130C12F412DC12C412AC1294",
		INIT_0D => X"1578156115491531151A150214EA14D214BB14A3148B1473145B1443142C1414",
		INIT_0E => X"16F216DA16C316AB1694167C1665164D1635161E160615EF15D715BF15A81590",
		INIT_0F => X"1867185018391821180A17F317DC17C417AD1795177E1767174F173817201709",
		INIT_10 => X"19D919C219AB1994197D1966194F19381921190A18F218DB18C418AD1896187E",
		INIT_11 => X"1B471B301B191B031AEC1AD51ABE1AA71A911A7A1A631A4C1A351A1E1A0719F0",
		INIT_12 => X"1CB11C9A1C841C6D1C571C401C2A1C131BFC1BE61BCF1BB81BA21B8B1B741B5E",
		INIT_13 => X"1E161E001DEA1DD31DBD1DA71D911D7A1D641D4E1D371D211D0A1CF41CDE1CC7",
		INIT_14 => X"1F771F611F4B1F351F1F1F091EF31EDD1EC71EB11E9B1E851E6F1E581E421E2C",
		INIT_15 => X"20D220BD20A72092207C20662050203B2025200F1FFA1FE41FCE1FB81FA21F8C",
		INIT_16 => X"2229221421FE21E921D421BE21A92194217E21692153213E2128211320FD20E8",
		INIT_17 => X"237A23662351233C2327231222FD22E722D222BD22A82293227E22692253223E",
		INIT_18 => X"24C624B2249D24892474245F244B24362421240C23F823E323CE23B923A4238F",
		INIT_19 => X"260D25F825E425D025BC25A72593257F256A25562541252D2519250424F024DB",
		INIT_1A => X"274D27392725271126FE26EA26D626C226AE269A26862671265D264926352621",
		INIT_1B => X"288728742860284D28392826281227FF27EB27D727C427B0279C278927752761",
		INIT_1C => X"29BC29A829952982296F295C294929362922290F28FC28E828D528C228AE289B",
		INIT_1D => X"2AE92AD72AC42AB12A9E2A8C2A792A662A532A402A2D2A1B2A0829F529E229CF",
		INIT_1E => X"2C102BFE2BEC2BD92BC72BB52BA22B902B7E2B6B2B592B462B342B212B0E2AFC",
		INIT_1F => X"2D302D1F2D0D2CFB2CE92CD72CC52CB32CA12C8F2C7D2C6B2C592C472C352C22",
		INIT_20 => X"2E4A2E382E272E162E042DF32DE12DD02DBE2DAC2D9B2D892D772D662D542D42",
		INIT_21 => X"2F5C2F4B2F3A2F292F182F072EF62EE52ED42EC32EB12EA02E8F2E7E2E6C2E5B",
		INIT_22 => X"30673056304630353025301430032FF32FE22FD12FC12FB02F9F2F8E2F7E2F6D",
		INIT_23 => X"316A315A314A313A312A311A310A30F930E930D930C930B930A8309830873077",
		INIT_24 => X"326632563247323732283218320831F931E931D931C931BA31AA319A318A317A",
		INIT_25 => X"335A334B333C332D331D330E32FF32F032E132D132C232B332A3329432853275",
		INIT_26 => X"344634373429341A340B33FD33EE33DF33D133C233B333A43395338733783369",
		INIT_27 => X"352A351C350E350034F134E334D534C734B934AA349C348E347F347134633454",
		INIT_28 => X"360535F835EA35DD35CF35C235B435A63599358B357D356F3561355435463538",
		INIT_29 => X"36D936CC36BF36B236A53698368B367D3670366336563648363B362E36203613",
		INIT_2A => X"37A43797378B377E377237653759374C373F373337263719370C370036F336E6",
		INIT_2B => X"3866385A384E38423836382A381E3812380637FA37EE37E137D537C937BD37B0",
		INIT_2C => X"39203915390938FE38F238E738DB38D038C438B938AD38A13895388A387E3872",
		INIT_2D => X"39D139C639BB39B039A5399A398F39843979396E39633958394D39423936392B",
		INIT_2E => X"3A793A6E3A643A5A3A503A453A3B3A303A263A1B3A113A0639FC39F139E639DB",
		INIT_2F => X"3B183B0E3B043AFA3AF13AE73ADD3AD33AC93ABF3AB53AAB3AA13A973A8D3A83",
		INIT_30 => X"3BAD3BA43B9B3B923B893B803B763B6D3B643B5A3B513B473B3E3B343B2B3B21",
		INIT_31 => X"3C3A3C313C293C203C183C0F3C063BFE3BF53BEC3BE33BDA3BD13BC83BBF3BB6",
		INIT_32 => X"3CBD3CB53CAD3CA53C9D3C953C8D3C853C7D3C753C6C3C643C5C3C533C4B3C42",
		INIT_33 => X"3D373D303D293D213D1A3D123D0B3D033CFB3CF43CEC3CE43CDD3CD53CCD3CC5",
		INIT_34 => X"3DA83DA13D9A3D933D8C3D863D7F3D783D713D6A3D633D5B3D543D4D3D463D3F",
		INIT_35 => X"3E0F3E093E023DFC3DF63DF03DE93DE33DDC3DD63DCF3DC93DC23DBC3DB53DAE",
		INIT_36 => X"3E6C3E673E613E5B3E563E503E4A3E443E3F3E393E333E2D3E273E213E1B3E15",
		INIT_37 => X"3EC03EBB3EB63EB13EAC3EA73EA23E9C3E973E923E8D3E873E823E7D3E773E72",
		INIT_38 => X"3F0A3F063F013EFD3EF83EF43EEF3EEB3EE63EE13EDD3ED83ED33ECE3ECA3EC5",
		INIT_39 => X"3F4A3F473F433F3F3F3B3F373F333F2F3F2B3F273F233F1F3F1B3F173F133F0E",
		INIT_3A => X"3F813F7E3F7B3F773F743F713F6E3F6A3F673F633F603F5C3F593F553F523F4E",
		INIT_3B => X"3FAE3FAB3FA93FA63FA33FA13F9E3F9B3F993F963F933F903F8D3F8A3F873F84",
		INIT_3C => X"3FD13FCF3FCD3FCB3FC93FC73FC53FC33FC03FBE3FBC3FBA3FB73FB53FB33FB0",
		INIT_3D => X"3FEA3FE93FE73FE63FE43FE33FE23FE03FDE3FDD3FDB3FDA3FD83FD63FD43FD3",
		INIT_3E => X"3FF93FF83FF83FF73FF63FF53FF53FF43FF33FF23FF13FF03FEF3FED3FEC3FEB",
		INIT_3F => X"3FFE3FFE3FFE3FFE3FFE3FFE3FFE3FFD3FFD3FFD3FFC3FFC3FFB3FFB3FFA3FFA",

      -- INIT_A/INIT_B: Initial values on output port
      INIT_A => X"000000000",
      INIT_B => X"000000000",
      -- INIT_FILE: Optional file used to specify initial RAM contents
      INIT_FILE => "NONE",
      -- RSTTYPE: "SYNC" or "ASYNC" 
      RSTTYPE => "SYNC",
      -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
      RST_PRIORITY_A => "CE",
      RST_PRIORITY_B => "CE",
      -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
      SIM_COLLISION_CHECK => "ALL",
      -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
      SIM_DEVICE => "SPARTAN6",
      -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
      SRVAL_A => X"000000000",
      SRVAL_B => X"000000000",
      -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
      WRITE_MODE_A => "READ_FIRST",
      WRITE_MODE_B => "READ_FIRST" 
   )
   port map (
      -- Port A Data: 32-bit (each) output: Port A data
      DOA => DOA_OUT,       -- 32-bit output: A port data output
      DOPA => DOPA_OUT,     -- 4-bit output: A port parity output
      -- Port B Data: 32-bit (each) output: Port B data
      DOB => DOB,       -- 32-bit output: B port data output
      DOPB => DOPB,     -- 4-bit output: B port parity output
      -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
      ADDRA => ADDRA_IN,   -- 14-bit input: A port address input
      CLKA => CLK_IN,     -- 1-bit input: A port clock input
      ENA => ENA_IN,       -- 1-bit input: A port enable input
      REGCEA => REGCEA, -- 1-bit input: A port register clock enable input
      RSTA => RSTA,     -- 1-bit input: A port register set/reset input
      WEA => WEA,       -- 4-bit input: Port A byte-wide write enable input
      -- Port A Data: 32-bit (each) input: Port A data
      DIA => DIA,       -- 32-bit input: A port data input
      DIPA => DIPA,     -- 4-bit input: A port parity input
      -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
      ADDRB => ADDRB_IN,   -- 14-bit input: B port address input
      CLKB => CLK_IN,     -- 1-bit input: B port clock input
      ENB => ENB_IN,       -- 1-bit input: B port enable input
      REGCEB => REGCEB, -- 1-bit input: B port register clock enable input
      RSTB => RSTB,     -- 1-bit input: B port register set/reset input
      WEB => WEB,       -- 4-bit input: Port B byte-wide write enable input
      -- Port B Data: 32-bit (each) input: Port B data
      DIB => DIB_IN,       -- 32-bit input: B port data input
      DIPB => DIPB_IN      -- 4-bit input: B port parity input
   );


   -- End of RAMB16BWER_inst instantiation
end Behavioral;

