----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:07:53 11/05/2021 
-- Design Name: 
-- Module Name:    BRAMHandler - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity BRAMHandler_CurveA_B01 is
	 Generic ( DataWidth : integer := 18);
    Port ( CLK_IN : in  STD_LOGIC;
			  ENA_IN : in STD_LOGIC;
           ADDRA_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DOA_OUT : out  STD_LOGIC_VECTOR(31 downto 0);
			  DOPA_OUT : out  STD_LOGIC_VECTOR(3 downto 0);
			  ENB_IN : in STD_LOGIC;
           ADDRB_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DIB_IN : in  STD_LOGIC_VECTOR(31 downto 0);
			  DIPB_IN : in  STD_LOGIC_VECTOR(3 downto 0));
end BRAMHandler_CurveA_B01;

architecture Behavioral of BRAMHandler_CurveA_B01 is

	signal REGCEA: STD_LOGIC := '0';
	signal RSTA: STD_LOGIC := '0';
	signal WEA : STD_LOGIC_VECTOR(3 downto 0)  := (others => '0');
	signal DIA : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DIPA : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');

	signal DOB : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DOPB : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');
	signal REGCEB: STD_LOGIC := '0';
	signal RSTB: STD_LOGIC := '0';
	signal WEB : STD_LOGIC_VECTOR(3 downto 0) := (others => '1');
	
begin

	-- RAMB16BWER: 16k-bit Data and 2k-bit Parity Configurable Synchronous Dual Port Block RAM with Optional Output Registers
   --             Spartan-6
   -- Xilinx HDL Language Template, version 14.7

   RAMB16BWER_inst01 : RAMB16BWER
   generic map (
      -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
      DATA_WIDTH_A => DataWidth,
      DATA_WIDTH_B => DataWidth,
      -- DOA_REG/DOB_REG: Optional output register (0 or 1)
      DOA_REG => 0,
      DOB_REG => 0,
      -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
      EN_RSTRAM_A => TRUE,
      EN_RSTRAM_B => TRUE,
     	-- INITP_00 to INITP_07: Initial memory contents.
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

		-- INIT_00 to INIT_3F: Initial memory contents.
		INIT_00 => X"7FF67FF77FF87FF97FFA7FFA7FFB7FFC7FFC7FFD7FFD7FFE7FFE7FFE7FFE7FFE",
		INIT_01 => X"7FD97FDB7FDE7FE07FE27FE47FE67FE87FEA7FEB7FED7FEF7FF07FF27FF37FF4",
		INIT_02 => X"7FA87FAC7FB07FB37FB67FBA7FBD7FC07FC37FC67FC97FCC7FCF7FD17FD47FD6",
		INIT_03 => X"7F647F697F6E7F737F777F7C7F807F857F897F8D7F917F957F997F9D7FA17FA5",
		INIT_04 => X"7F0D7F137F197F1F7F247F2A7F307F357F3B7F407F467F4B7F507F557F5A7F5F",
		INIT_05 => X"7EA17EA87EB07EB77EBE7EC57ECC7ED37ED97EE07EE77EED7EF47EFA7F007F06",
		INIT_06 => X"7E227E2B7E337E3C7E447E4C7E547E5C7E647E6C7E747E7C7E837E8B7E927E9A",
		INIT_07 => X"7D907D9A7DA37DAD7DB67DC07DC97DD27DDC7DE57DEE7DF77E007E087E117E1A",
		INIT_08 => X"7CEA7CF57D007D0B7D157D207D2B7D357D3F7D4A7D547D5E7D687D727D7C7D86",
		INIT_09 => X"7C317C3D7C497C557C617C6D7C797C847C907C9C7CA77CB27CBE7CC97CD47CDF",
		INIT_0A => X"7B657B727B807B8D7B9A7BA77BB47BC17BCD7BDA7BE77BF37C007C0C7C197C25",
		INIT_0B => X"7A867A947AA37AB17ABF7ACE7ADC7AEA7AF87B067B147B217B2F7B3D7B4A7B58",
		INIT_0C => X"799479A379B379C379D279E179F17A007A0F7A1E7A2D7A3C7A4B7A5A7A697A77",
		INIT_0D => X"788F78A078B078C178D278E278F3790379147924793479447954796479747984",
		INIT_0E => X"77777789779B77AD77BF77D177E277F47805781778287839784B785C786D787E",
		INIT_0F => X"764D766176747687769A76AD76BF76D276E576F7770A771C772F774177537765",
		INIT_10 => X"75117526753A754E75627576758A759E75B275C575D975ED760076147627763A",
		INIT_11 => X"73C373D973EE74037418742D74437458746C7481749674AB74BF74D474E974FD",
		INIT_12 => X"7263727A729072A672BD72D372E972FF7315732B73417357736D7382739873AE",
		INIT_13 => X"70F1710971207138714F7167717E719571AC71C371DA71F17208721F7236724C",
		INIT_14 => X"6F6E6F876FA06FB86FD16FE97001701A7032704A7062707A709270AA70C270DA",
		INIT_15 => X"6DDA6DF46E0D6E276E416E5A6E736E8D6EA66EBF6ED96EF26F0B6F246F3D6F55",
		INIT_16 => X"6C356C4F6C6A6C856C9F6CBA6CD56CEF6D096D246D3E6D586D726D8C6DA66DC0",
		INIT_17 => X"6A7F6A9A6AB66AD26AEE6B096B256B406B5C6B776B926BAD6BC96BE46BFF6C1A",
		INIT_18 => X"68B868D568F2690F692B694869646981699D69BA69D669F26A0F6A2B6A476A63",
		INIT_19 => X"66E266FF671D673B67596776679467B167CF67EC680A682768446861687E689B",
		INIT_1A => X"64FB651A653965586576659565B365D265F0660F662D664B6669668866A666C4",
		INIT_1B => X"6305632563456364638463A463C363E36402642164416460647F649E64BD64DC",
		INIT_1C => X"6100612161416162618361A361C461E46204622562456265628562A562C562E5",
		INIT_1D => X"5EEC5F0D5F2F5F515F725F945FB55FD65FF86019603A605B607C609D60BE60DF",
		INIT_1E => X"5CC95CEB5D0E5D305D535D755D975DBA5DDC5DFE5E205E425E645E865EA85ECA",
		INIT_1F => X"5A975ABB5ADE5B025B255B485B6C5B8F5BB25BD55BF85C1B5C3E5C615C835CA6",
		INIT_20 => X"5858587D58A158C558E9590E59325956597A599E59C159E55A095A2D5A505A74",
		INIT_21 => X"560B56315656567B56A056C556EA570F57345758577D57A257C657EB580F5834",
		INIT_22 => X"53B153D753FD54235449546F549554BA54E05506552B55515576559C55C155E6",
		INIT_23 => X"514A5171519851BF51E5520C52325259527F52A652CC52F35319533F5365538B",
		INIT_24 => X"4ED74EFE4F264F4D4F754F9C4FC44FEB501250395060508850AF50D650FD5123",
		INIT_25 => X"4C574C7F4CA84CD04CF84D204D484D704D984DC04DE84E104E384E604E874EAF",
		INIT_26 => X"49CC49F54A1E4A474A704A984AC14AEA4B134B3B4B644B8D4BB54BDE4C064C2F",
		INIT_27 => X"4735475E478847B247DB4805482F4858488248AB48D448FE49274950497949A2",
		INIT_28 => X"449344BD44E84512453C4567459145BB45E5460F46394663468D46B746E1470B",
		INIT_29 => X"41E64211423C4267429242BD42E84313433E4369439343BE43E94413443E4468",
		INIT_2A => X"3F303F5B3F873FB33FDE400A40354061408C40B840E3410E413A4165419041BB",
		INIT_2B => X"3C6F3C9C3CC83CF43D203D4D3D793DA53DD13DFD3E293E553E813EAC3ED83F04",
		INIT_2C => X"39A639D339FF3A2C3A593A863AB23ADF3B0C3B383B653B913BBE3BEA3C173C43",
		INIT_2D => X"36D33701372E375B378937B637E33810383D386B389838C538F2391F394C3979",
		INIT_2E => X"33F834263454348234B034DD350B35393567359435C235F0361D364B367836A6",
		INIT_2F => X"31153143317231A031CF31FD322B3259328832B632E433123340336E339C33CA",
		INIT_30 => X"2E2A2E592E882EB72EE62F142F432F722FA12FCF2FFE302C305B308A30B830E7",
		INIT_31 => X"2B392B682B972BC62BF62C252C542C832CB22CE12D112D402D6F2D9E2DCD2DFB",
		INIT_32 => X"2840287028A028CF28FF292F295E298E29BD29ED2A1C2A4C2A7B2AAB2ADA2B09",
		INIT_33 => X"2542257225A225D2260226322662269226C226F227212751278127B127E12810",
		INIT_34 => X"223D226E229E22CE22FF232F235F239023C023F024212451248124B124E12511",
		INIT_35 => X"1F341F641F951FC61FF620272058208820B920EA211A214B217B21AC21DC220D",
		INIT_36 => X"1C251C561C871CB81CE91D1A1D4B1D7C1DAD1DDE1E0F1E3F1E701EA11ED21F03",
		INIT_37 => X"19121944197519A619D71A091A3A1A6B1A9C1ACD1AFE1B301B611B921BC31BF4",
		INIT_38 => X"15FC162D165F169016C216F317241756178717B917EA181C184D187E18B018E1",
		INIT_39 => X"12E113131345137713A813DA140C143D146F14A114D2150415351567159815CA",
		INIT_3A => X"0FC40FF61028105A108C10BE10F011211153118511B711E9121A124C127E12B0",
		INIT_3B => X"0CA50CD70D090D3B0D6D0D9F0DD10E030E350E670E990ECB0EFD0F2F0F610F93",
		INIT_3C => X"098409B609E80A1A0A4C0A7E0AB00AE20B150B470B790BAB0BDD0C0F0C410C73",
		INIT_3D => X"0661069306C506F7072A075C078E07C007F208250857088908BB08ED091F0952",
		INIT_3E => X"033D036F03A103D404060438046A049D04CF050105330566059805CA05FC062F",
		INIT_3F => X"0019004B007D00AF00E201140146017901AB01DD020F0242027402A602D8030B",
      -- INIT_A/INIT_B: Initial values on output port
      INIT_A => X"000000000",
      INIT_B => X"000000000",
      -- INIT_FILE: Optional file used to specify initial RAM contents
      INIT_FILE => "NONE",
      -- RSTTYPE: "SYNC" or "ASYNC" 
      RSTTYPE => "SYNC",
      -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
      RST_PRIORITY_A => "CE",
      RST_PRIORITY_B => "CE",
      -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
      SIM_COLLISION_CHECK => "ALL",
      -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
      SIM_DEVICE => "SPARTAN6",
      -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
      SRVAL_A => X"000000000",
      SRVAL_B => X"000000000",
      -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
      WRITE_MODE_A => "READ_FIRST",
      WRITE_MODE_B => "READ_FIRST" 
   )
   port map (
      -- Port A Data: 32-bit (each) output: Port A data
      DOA => DOA_OUT,       -- 32-bit output: A port data output
      DOPA => DOPA_OUT,     -- 4-bit output: A port parity output
      -- Port B Data: 32-bit (each) output: Port B data
      DOB => DOB,       -- 32-bit output: B port data output
      DOPB => DOPB,     -- 4-bit output: B port parity output
      -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
      ADDRA => ADDRA_IN,   -- 14-bit input: A port address input
      CLKA => CLK_IN,     -- 1-bit input: A port clock input
      ENA => ENA_IN,       -- 1-bit input: A port enable input
      REGCEA => REGCEA, -- 1-bit input: A port register clock enable input
      RSTA => RSTA,     -- 1-bit input: A port register set/reset input
      WEA => WEA,       -- 4-bit input: Port A byte-wide write enable input
      -- Port A Data: 32-bit (each) input: Port A data
      DIA => DIA,       -- 32-bit input: A port data input
      DIPA => DIPA,     -- 4-bit input: A port parity input
      -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
      ADDRB => ADDRB_IN,   -- 14-bit input: B port address input
      CLKB => CLK_IN,     -- 1-bit input: B port clock input
      ENB => ENB_IN,       -- 1-bit input: B port enable input
      REGCEB => REGCEB, -- 1-bit input: B port register clock enable input
      RSTB => RSTB,     -- 1-bit input: B port register set/reset input
      WEB => WEB,       -- 4-bit input: Port B byte-wide write enable input
      -- Port B Data: 32-bit (each) input: Port B data
      DIB => DIB_IN,       -- 32-bit input: B port data input
      DIPB => DIPB_IN      -- 4-bit input: B port parity input
   );

   -- End of RAMB16BWER_inst instantiation
end Behavioral;

