----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:07:53 11/05/2021 
-- Design Name: 
-- Module Name:    BRAMHandler - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity BRAMHandler_CurveA_B11 is
	 Generic ( DataWidth : integer := 18);
    Port ( CLK_IN : in  STD_LOGIC;
			  ENA_IN : in STD_LOGIC;
           ADDRA_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DOA_OUT : out  STD_LOGIC_VECTOR(31 downto 0);
			  DOPA_OUT : out  STD_LOGIC_VECTOR(3 downto 0);
			  ENB_IN : in STD_LOGIC;
           ADDRB_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DIB_IN : in  STD_LOGIC_VECTOR(31 downto 0);
			  DIPB_IN : in  STD_LOGIC_VECTOR(3 downto 0));
end BRAMHandler_CurveA_B11;

architecture Behavioral of BRAMHandler_CurveA_B11 is

	signal REGCEA: STD_LOGIC := '0';
	signal RSTA: STD_LOGIC := '0';
	signal WEA : STD_LOGIC_VECTOR(3 downto 0)  := (others => '0');
	signal DIA : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DIPA : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');

	signal DOB : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DOPB : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');
	signal REGCEB: STD_LOGIC := '0';
	signal RSTB: STD_LOGIC := '0';
	signal WEB : STD_LOGIC_VECTOR(3 downto 0) := (others => '1');
	
begin

	-- RAMB16BWER: 16k-bit Data and 2k-bit Parity Configurable Synchronous Dual Port Block RAM with Optional Output Registers
   --             Spartan-6
   -- Xilinx HDL Language Template, version 14.7

   RAMB16BWER_inst11 : RAMB16BWER
   generic map (
      -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
      DATA_WIDTH_A => DataWidth,
      DATA_WIDTH_B => DataWidth,
      -- DOA_REG/DOB_REG: Optional output register (0 or 1)
      DOA_REG => 0,
      DOB_REG => 0,
      -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
      EN_RSTRAM_A => TRUE,
      EN_RSTRAM_B => TRUE,
      -- INITP_00 to INITP_07: Initial memory contents.
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

		-- INIT_00 to INIT_3F: Initial memory contents.
		INIT_00 => X"800B800A80098008800780068005800480048003800380028002800280028002",
		INIT_01 => X"8028802680248021801F801D801B801980178015801480128011800F800E800C",
		INIT_02 => X"805980568052804F804B804880458042803E803B8038803680338030802D802B",
		INIT_03 => X"809E809980948090808B80878082807E807980758071806D806980658061805D",
		INIT_04 => X"80F780F080EA80E480DF80D980D380CD80C880C280BD80B880B280AD80A880A3",
		INIT_05 => X"8162815B8154814D8146813F81388131812A8123811D811681108109810380FD",
		INIT_06 => X"81E281D981D181C981C081B881B081A881A0819881908188818181798171816A",
		INIT_07 => X"8275826B82628258824E8245823C8232822982208217820E820581FC81F381EB",
		INIT_08 => X"831B8310830582FB82F082E582DB82D082C682BB82B182A7829D82938289827F",
		INIT_09 => X"83D583C983BD83B183A58399838D83818376836A835F83538348833D83318326",
		INIT_0A => X"84A284948487847A846D8460845384468439842C841F8413840683FA83ED83E1",
		INIT_0B => X"858185738564855685488539852B851D850F850184F384E684D884CA84BD84AF",
		INIT_0C => X"8674866486558645863686268617860885F885E985DA85CB85BC85AE859F8590",
		INIT_0D => X"877A876987588747873787268715870586F586E486D486C486B486A486948684",
		INIT_0E => X"88928880886E885C884A883888268815880387F287E087CF87BE87AD879C878B",
		INIT_0F => X"89BC89A9899689838970895D894A89378925891288FF88ED88DB88C888B688A4",
		INIT_10 => X"8AF98AE58AD08ABC8AA88A948A808A6C8A588A448A318A1D8A0A89F689E389CF",
		INIT_11 => X"8C488C328C1D8C078BF28BDD8BC88BB38B9E8B898B748B608B4B8B368B228B0D",
		INIT_12 => X"8DA88D928D7B8D658D4E8D388D228D0C8CF68CE08CCA8CB48C9E8C888C738C5D",
		INIT_13 => X"8F1B8F038EEB8ED48EBC8EA58E8E8E768E5F8E488E318E1A8E038DEC8DD68DBF",
		INIT_14 => X"909E9085906D9054903C9023900B8FF28FDA8FC28FAA8F928F7A8F628F4A8F32",
		INIT_15 => X"92339219920091E691CC91B3919991809166914D9134911B910290E990D090B7",
		INIT_16 => X"93D993BE93A39389936E93539339931E930492EA92CF92B5929B92819267924D",
		INIT_17 => X"958F95739558953C9520950594E994CD94B29497947B94609445942A940F93F4",
		INIT_18 => X"97569739971D970096E396C696AA968D967196549638961C960095E395C795AB",
		INIT_19 => X"992D990F98F298D498B69898987B985D98409822980597E897CB97AD97909773",
		INIT_1A => X"9B149AF59AD79AB89A999A7A9A5C9A3D9A1F9A0099E299C499A699879969994B",
		INIT_1B => X"9D0B9CEB9CCB9CAB9C8C9C6C9C4D9C2D9C0E9BEE9BCF9BB09B909B719B529B33",
		INIT_1C => X"9F119EF09ECF9EAE9E8E9E6D9E4D9E2C9E0C9DEB9DCB9DAB9D8B9D6B9D4B9D2B",
		INIT_1D => X"A125A104A0E2A0C0A09FA07DA05CA03AA0199FF89FD79FB59F949F739F529F31",
		INIT_1E => X"A349A326A303A2E1A2BEA29CA27AA257A235A213A1F1A1CFA1ADA18BA169A147",
		INIT_1F => X"A57AA557A533A510A4EDA4C9A4A6A483A460A43DA41AA3F7A3D4A3B1A38EA36B",
		INIT_20 => X"A7BAA796A771A74DA729A705A6E0A6BCA698A674A651A62DA609A5E5A5C1A59E",
		INIT_21 => X"AA07A9E2A9BDA998A973A94EA929A904A8DFA8BAA895A871A84CA827A803A7DE",
		INIT_22 => X"AC62AC3CAC16ABF0ABCAABA4AB7EAB58AB33AB0DAAE8AAC2AA9DAA77AA52AA2C",
		INIT_23 => X"AEC9AEA2AE7BAE55AE2EAE07ADE1ADBAAD94AD6DAD47AD21ACFAACD4ACAEAC88",
		INIT_24 => X"B13DB115B0EEB0C6B09FB077B050B029B002AFDAAFB3AF8CAF65AF3EAF17AEF0",
		INIT_25 => X"B3BDB395B36CB344B31CB2F4B2CCB2A4B27CB254B22CB204B1DCB1B4B18CB165",
		INIT_26 => X"B649B620B5F7B5CEB5A5B57CB553B52AB502B4D9B4B0B488B45FB436B40EB3E6",
		INIT_27 => X"B8E0B8B6B88DB863B839B810B7E6B7BDB793B76AB740B717B6EEB6C4B69BB672",
		INIT_28 => X"BB82BB58BB2EBB03BAD9BAAFBA84BA5ABA30BA06B9DCB9B2B988B95EB934B90A",
		INIT_29 => X"BE2FBE04BDD9BDAEBD83BD58BD2DBD02BCD8BCADBC82BC57BC2DBC02BBD7BBAD",
		INIT_2A => X"C0E6C0BAC08FC063C037C00CBFE0BFB5BF89BF5EBF33BF07BEDCBEB1BE86BE5A",
		INIT_2B => X"C3A7C37AC34EC322C2F6C2CAC29DC271C245C219C1EDC1C1C195C16AC13EC112",
		INIT_2C => X"C671C644C617C5EAC5BDC591C564C537C50BC4DEC4B1C485C458C42CC400C3D3",
		INIT_2D => X"C944C916C8E9C8BBC88EC861C834C806C7D9C7ACC77FC752C725C6F8C6CBC69E",
		INIT_2E => X"CC1FCBF1CBC3CB95CB67CB39CB0CCADECAB0CA83CA55CA27C9FAC9CCC99FC971",
		INIT_2F => X"CF02CED4CEA5CE77CE49CE1ACDECCDBECD90CD61CD33CD05CCD7CCA9CC7BCC4D",
		INIT_30 => X"D1EDD1BED18FD160D132D103D0D4D0A5D077D048D019CFEBCFBCCF8ECF5FCF31",
		INIT_31 => X"D4DFD4B0D480D451D422D3F3D3C3D394D365D336D307D2D8D2A9D27AD24BD21C",
		INIT_32 => X"D7D8D7A8D778D749D719D6E9D6BAD68AD65BD62BD5FCD5CCD59DD56DD53ED50E",
		INIT_33 => X"DAD6DAA6DA76DA46DA16D9E6D9B6D986D956D926D8F7D8C7D897D867D837D807",
		INIT_34 => X"DDDBDDABDD7ADD4ADD19DCE9DCB9DC88DC58DC28DBF8DBC7DB97DB67DB37DB07",
		INIT_35 => X"E0E5E0B4E083E053E022DFF1DFC1DF90DF5FDF2FDEFEDECEDE9DDE6CDE3CDE0C",
		INIT_36 => X"E3F3E3C2E391E360E32FE2FEE2CDE29DE26CE23BE20AE1D9E1A8E177E146E116",
		INIT_37 => X"E706E6D5E6A4E673E641E610E5DFE5AEE57CE54BE51AE4E9E4B8E487E456E425",
		INIT_38 => X"EA1DE9ECE9BAE989E957E926E8F4E8C3E891E860E82FE7FDE7CCE79AE769E738",
		INIT_39 => X"ED37ED06ECD4ECA2EC71EC3FEC0DEBDCEBAAEB78EB47EB15EAE3EAB2EA80EA4F",
		INIT_3A => X"F054F023EFF1EFBFEF8DEF5BEF29EEF7EEC6EE94EE62EE30EDFEEDCDED9BED69",
		INIT_3B => X"F374F342F310F2DEF2ACF27AF248F216F1E4F1B2F180F14EF11CF0EAF0B8F086",
		INIT_3C => X"F695F663F631F5FFF5CDF59BF569F537F504F4D2F4A0F46EF43CF40AF3D8F3A6",
		INIT_3D => X"F9B8F986F954F922F8EFF8BDF88BF859F827F7F5F7C2F790F75EF72CF6FAF6C8",
		INIT_3E => X"FCDCFCAAFC78FC45FC13FBE1FBAFFB7CFB4AFB18FAE6FAB3FA81FA4FFA1DF9EB",
		INIT_3F => X"0000FFCEFF9CFF6AFF37FF05FED3FEA1FE6EFE3CFE0AFDD7FDA5FD73FD41FD0E",
      -- INIT_A/INIT_B: Initial values on output port
      INIT_A => X"000000000",
      INIT_B => X"000000000",
      -- INIT_FILE: Optional file used to specify initial RAM contents
      INIT_FILE => "NONE",
      -- RSTTYPE: "SYNC" or "ASYNC" 
      RSTTYPE => "SYNC",
      -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
      RST_PRIORITY_A => "CE",
      RST_PRIORITY_B => "CE",
      -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
      SIM_COLLISION_CHECK => "ALL",
      -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
      SIM_DEVICE => "SPARTAN6",
      -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
      SRVAL_A => X"000000000",
      SRVAL_B => X"000000000",
      -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
      WRITE_MODE_A => "READ_FIRST",
      WRITE_MODE_B => "READ_FIRST" 
   )
   port map (
      -- Port A Data: 32-bit (each) output: Port A data
      DOA => DOA_OUT,       -- 32-bit output: A port data output
      DOPA => DOPA_OUT,     -- 4-bit output: A port parity output
      -- Port B Data: 32-bit (each) output: Port B data
      DOB => DOB,       -- 32-bit output: B port data output
      DOPB => DOPB,     -- 4-bit output: B port parity output
      -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
      ADDRA => ADDRA_IN,   -- 14-bit input: A port address input
      CLKA => CLK_IN,     -- 1-bit input: A port clock input
      ENA => ENA_IN,       -- 1-bit input: A port enable input
      REGCEA => REGCEA, -- 1-bit input: A port register clock enable input
      RSTA => RSTA,     -- 1-bit input: A port register set/reset input
      WEA => WEA,       -- 4-bit input: Port A byte-wide write enable input
      -- Port A Data: 32-bit (each) input: Port A data
      DIA => DIA,       -- 32-bit input: A port data input
      DIPA => DIPA,     -- 4-bit input: A port parity input
      -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
      ADDRB => ADDRB_IN,   -- 14-bit input: B port address input
      CLKB => CLK_IN,     -- 1-bit input: B port clock input
      ENB => ENB_IN,       -- 1-bit input: B port enable input
      REGCEB => REGCEB, -- 1-bit input: B port register clock enable input
      RSTB => RSTB,     -- 1-bit input: B port register set/reset input
      WEB => WEB,       -- 4-bit input: Port B byte-wide write enable input
      -- Port B Data: 32-bit (each) input: Port B data
      DIB => DIB_IN,       -- 32-bit input: B port data input
      DIPB => DIPB_IN      -- 4-bit input: B port parity input
   );

   -- End of RAMB16BWER_inst instantiation
end Behavioral;

