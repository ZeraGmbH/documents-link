----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:07:53 11/05/2021 
-- Design Name: 
-- Module Name:    BRAMHandler - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity BRAMHandler_CurveA_B10 is
	 Generic ( DataWidth : integer := 18);
    Port ( CLK_IN : in  STD_LOGIC;
			  ENA_IN : in STD_LOGIC;
           ADDRA_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DOA_OUT : out  STD_LOGIC_VECTOR(31 downto 0);
			  DOPA_OUT : out  STD_LOGIC_VECTOR(3 downto 0);
			  ENB_IN : in STD_LOGIC;
           ADDRB_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DIB_IN : in  STD_LOGIC_VECTOR(31 downto 0);
			  DIPB_IN : in  STD_LOGIC_VECTOR(3 downto 0));
end BRAMHandler_CurveA_B10;

architecture Behavioral of BRAMHandler_CurveA_B10 is

	signal REGCEA: STD_LOGIC := '0';
	signal RSTA: STD_LOGIC := '0';
	signal WEA : STD_LOGIC_VECTOR(3 downto 0)  := (others => '0');
	signal DIA : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DIPA : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');

	signal DOB : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DOPB : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');
	signal REGCEB: STD_LOGIC := '0';
	signal RSTB: STD_LOGIC := '0';
	signal WEB : STD_LOGIC_VECTOR(3 downto 0) := (others => '1');
	
begin

	-- RAMB16BWER: 16k-bit Data and 2k-bit Parity Configurable Synchronous Dual Port Block RAM with Optional Output Registers
   --             Spartan-6
   -- Xilinx HDL Language Template, version 14.7

   RAMB16BWER_inst10 : RAMB16BWER
   generic map (
      -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
      DATA_WIDTH_A => DataWidth,
      DATA_WIDTH_B => DataWidth,
      -- DOA_REG/DOB_REG: Optional output register (0 or 1)
      DOA_REG => 0,
      DOB_REG => 0,
      -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
      EN_RSTRAM_A => TRUE,
      EN_RSTRAM_B => TRUE,
     	-- INITP_00 to INITP_07: Initial memory contents.
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

		-- INIT_00 to INIT_3F: Initial memory contents.
		INIT_00 => X"FCF5FD28FD5AFD8CFDBEFDF1FE23FE55FE87FEBAFEECFF1EFF51FF83FFB5FFE7",
		INIT_01 => X"F9D1FA04FA36FA68FA9AFACDFAFFFB31FB63FB96FBC8FBFAFC2CFC5FFC91FCC3",
		INIT_02 => X"F6AEF6E1F713F745F777F7A9F7DBF80EF840F872F8A4F8D6F909F93BF96DF99F",
		INIT_03 => X"F38DF3BFF3F1F423F455F487F4B9F4EBF51EF550F582F5B4F5E6F618F64AF67C",
		INIT_04 => X"F06DF09FF0D1F103F135F167F199F1CBF1FDF22FF261F293F2C5F2F7F329F35B",
		INIT_05 => X"ED50ED82EDB4EDE6EE17EE49EE7BEEADEEDFEF10EF42EF74EFA6EFD8F00AF03C",
		INIT_06 => X"EA36EA68EA99EACBEAFCEB2EEB5FEB91EBC3EBF4EC26EC58EC89ECBBECEDED1F",
		INIT_07 => X"E71FE750E782E7B3E7E4E816E847E879E8AAE8DCE90DE93EE970E9A1E9D3EA04",
		INIT_08 => X"E40CE43DE46EE49FE4D0E502E533E564E595E5C6E5F7E629E65AE68BE6BCE6EE",
		INIT_09 => X"E0FDE12EE15FE190E1C1E1F1E222E253E284E2B5E2E6E317E348E379E3AAE3DB",
		INIT_0A => X"DDF3DE24DE54DE85DEB5DEE6DF16DF47DF78DFA8DFD9E00AE03AE06BE09CE0CC",
		INIT_0B => X"DAEFDB1FDB4FDB7FDBAFDBDFDC10DC40DC70DCA1DCD1DD01DD32DD62DD92DDC3",
		INIT_0C => X"D7F0D81FD84FD87FD8AFD8DFD90ED93ED96ED99ED9CED9FEDA2EDA5EDA8EDABE",
		INIT_0D => X"D4F7D526D555D585D5B4D5E4D613D643D672D6A2D6D1D701D731D760D790D7C0",
		INIT_0E => X"D205D233D262D291D2C0D2EFD31FD34ED37DD3ACD3DBD40AD43AD469D498D4C7",
		INIT_0F => X"CF19CF48CF76CFA5CFD4D002D031D05FD08ED0BDD0ECD11AD149D178D1A7D1D6",
		INIT_10 => X"CC36CC64CC92CCC0CCEECD1CCD4ACD78CDA7CDD5CE03CE31CE60CE8ECEBDCEEB",
		INIT_11 => X"C95AC988C9B5C9E3CA10CA3ECA6CCA99CAC7CAF5CB23CB50CB7ECBACCBDACC08",
		INIT_12 => X"C687C6B4C6E1C70EC73BC768C795C7C3C7F0C81DC84AC877C8A5C8D2C8FFC92D",
		INIT_13 => X"C3BDC3E9C416C442C46FC49BC4C8C4F4C521C54EC57AC5A7C5D4C601C62DC65A",
		INIT_14 => X"C0FCC128C154C17FC1ABC1D7C203C22FC25BC287C2B3C2E0C30CC338C364C391",
		INIT_15 => X"BE45BE70BE9BBEC6BEF2BF1DBF48BF74BF9FBFCBBFF6C022C04DC079C0A5C0D0",
		INIT_16 => X"BB98BBC2BBEDBC17BC42BC6DBC97BCC2BCEDBD18BD43BD6EBD99BDC4BDEFBE1A",
		INIT_17 => X"B8F5B91FB949B973B99DB9C7B9F1BA1BBA45BA6FBA99BAC4BAEEBB18BB43BB6D",
		INIT_18 => X"B65EB687B6B0B6D9B702B72CB755B77EB7A8B7D1B7FBB825B84EB878B8A2B8CB",
		INIT_19 => X"B3D1B3FAB422B44BB473B49CB4C5B4EDB516B53FB568B590B5B9B5E2B60BB634",
		INIT_1A => X"B151B179B1A0B1C8B1F0B218B240B268B290B2B8B2E0B308B330B358B381B3A9",
		INIT_1B => X"AEDDAF03AF2AAF51AF78AFA0AFC7AFEEB015B03CB064B08BB0B3B0DAB102B129",
		INIT_1C => X"AC75AC9BACC1ACE7AD0DAD34AD5AAD81ADA7ADCEADF4AE1BAE41AE68AE8FAEB6",
		INIT_1D => X"AA1AAA3FAA64AA8AAAAFAAD5AAFAAB20AB46AB6BAB91ABB7ABDDAC03AC29AC4F",
		INIT_1E => X"A7CCA7F1A815A83AA85EA883A8A8A8CCA8F1A916A93BA960A985A9AAA9CFA9F5",
		INIT_1F => X"A58CA5B0A5D3A5F7A61BA63FA662A686A6AAA6CEA6F2A717A73BA75FA783A7A8",
		INIT_20 => X"A35AA37DA39FA3C2A3E5A408A42BA44EA471A494A4B8A4DBA4FEA522A545A569",
		INIT_21 => X"A136A158A17AA19CA1BEA1E0A202A224A246A269A28BA2ADA2D0A2F2A315A337",
		INIT_22 => X"9F219F429F639F849FA59FC69FE7A008A02AA04BA06CA08EA0AFA0D1A0F3A114",
		INIT_23 => X"9D1B9D3B9D5B9D7B9D9B9DBB9DDB9DFC9E1C9E3C9E5D9E7D9E9E9EBF9EDF9F00",
		INIT_24 => X"9B249B439B629B819BA09BBF9BDF9BFE9C1D9C3D9C5C9C7C9C9C9CBB9CDB9CFB",
		INIT_25 => X"993C995A9978999799B599D399F19A109A2E9A4D9A6B9A8A9AA89AC79AE69B05",
		INIT_26 => X"97659782979F97BC97D997F698149831984F986C988A98A798C598E39901991E",
		INIT_27 => X"959D95B995D595F1960E962A96469663967F969C96B896D596F1970E972B9748",
		INIT_28 => X"93E69401941C94379453946E948994A494C094DB94F79512952E954A95669581",
		INIT_29 => X"9240925A9274928E92A892C292DC92F79311932B93469361937B939693B193CB",
		INIT_2A => X"90AB90C390DC90F5910E91279141915A9173918D91A691BF91D991F3920C9226",
		INIT_2B => X"8F268F3E8F568F6E8F868F9E8FB68FCE8FE68FFF9017902F9048906090799092",
		INIT_2C => X"8DB48DCA8DE18DF88E0F8E268E3D8E548E6B8E828E998EB18EC88EE08EF78F0F",
		INIT_2D => X"8C528C688C7E8C938CA98CBF8CD58CEB8D018D178D2D8D438D5A8D708D868D9D",
		INIT_2E => X"8B038B178B2C8B418B558B6A8B7F8B948BA88BBD8BD38BE88BFD8C128C278C3D",
		INIT_2F => X"89C689D989EC8A008A138A278A3B8A4E8A628A768A8A8A9E8AB28AC68ADA8AEF",
		INIT_30 => X"889B88AD88BF88D188E488F68909891B892E8941895389668979898C899F89B3",
		INIT_31 => X"8782879387A487B587C787D887E987FB880C881E882F88418853886588778889",
		INIT_32 => X"867C868C869C86AC86BC86CC86DC86EC86FD870D871E872E873F875087608771",
		INIT_33 => X"8589859785A685B585C485D385E285F18600860F861F862E863D864D865D866C",
		INIT_34 => X"84A884B684C384D184DF84EC84FA85088516852485328541854F855D856C857A",
		INIT_35 => X"83DB83E783F48400840D841984268433843F844C8459846684738480848E849B",
		INIT_36 => X"8321832C83378342834E835983648370837C83878393839F83AB83B783C383CF",
		INIT_37 => X"827A8284828E829882A282AC82B682C182CB82D582E082EB82F58300830B8316",
		INIT_38 => X"81E681EF81F8820082098212821B8224822E82378240824A8253825D82668270",
		INIT_39 => X"8166816E8175817D8184818C8194819C81A481AC81B481BC81C481CD81D581DE",
		INIT_3A => X"80FA81008106810C8113811981208127812D8134813B8142814981508158815F",
		INIT_3B => X"80A180A680AB80B080B580BA80C080C580CB80D080D680DC80E180E780ED80F3",
		INIT_3C => X"805B805F80638067806B806F80738077807B808080848089808D80928097809C",
		INIT_3D => X"802A802C802F803180348037803A803D804080438046804A804D805080548058",
		INIT_3E => X"800C800D800E801080118013801580168018801A801C801E8020802280258027",
		INIT_3F => X"800280028002800280028003800380048004800580068006800780088009800A",
      -- INIT_A/INIT_B: Initial values on output port
      INIT_A => X"000000000",
      INIT_B => X"000000000",
      -- INIT_FILE: Optional file used to specify initial RAM contents
      INIT_FILE => "NONE",
      -- RSTTYPE: "SYNC" or "ASYNC" 
      RSTTYPE => "SYNC",
      -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
      RST_PRIORITY_A => "CE",
      RST_PRIORITY_B => "CE",
      -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
      SIM_COLLISION_CHECK => "ALL",
      -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
      SIM_DEVICE => "SPARTAN6",
      -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
      SRVAL_A => X"000000000",
      SRVAL_B => X"000000000",
      -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
      WRITE_MODE_A => "READ_FIRST",
      WRITE_MODE_B => "READ_FIRST" 
   )
   port map (
      -- Port A Data: 32-bit (each) output: Port A data
      DOA => DOA_OUT,       -- 32-bit output: A port data output
      DOPA => DOPA_OUT,     -- 4-bit output: A port parity output
      -- Port B Data: 32-bit (each) output: Port B data
      DOB => DOB,       -- 32-bit output: B port data output
      DOPB => DOPB,     -- 4-bit output: B port parity output
      -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
      ADDRA => ADDRA_IN,   -- 14-bit input: A port address input
      CLKA => CLK_IN,     -- 1-bit input: A port clock input
      ENA => ENA_IN,       -- 1-bit input: A port enable input
      REGCEA => REGCEA, -- 1-bit input: A port register clock enable input
      RSTA => RSTA,     -- 1-bit input: A port register set/reset input
      WEA => WEA,       -- 4-bit input: Port A byte-wide write enable input
      -- Port A Data: 32-bit (each) input: Port A data
      DIA => DIA,       -- 32-bit input: A port data input
      DIPA => DIPA,     -- 4-bit input: A port parity input
      -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
      ADDRB => ADDRB_IN,   -- 14-bit input: B port address input
      CLKB => CLK_IN,     -- 1-bit input: B port clock input
      ENB => ENB_IN,       -- 1-bit input: B port enable input
      REGCEB => REGCEB, -- 1-bit input: B port register clock enable input
      RSTB => RSTB,     -- 1-bit input: B port register set/reset input
      WEB => WEB,       -- 4-bit input: Port B byte-wide write enable input
      -- Port B Data: 32-bit (each) input: Port B data
      DIB => DIB_IN,       -- 32-bit input: B port data input
      DIPB => DIPB_IN      -- 4-bit input: B port parity input
   );

   -- End of RAMB16BWER_inst instantiation
end Behavioral;

