----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:07:53 11/05/2021 
-- Design Name: 
-- Module Name:    BRAMHandler - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity BRAMHandler_CurveA_B00 is
	 Generic ( DataWidth : integer := 18);
    Port ( CLK_IN : in  STD_LOGIC;
			  ENA_IN : in STD_LOGIC;
           ADDRA_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DOA_OUT : out  STD_LOGIC_VECTOR(31 downto 0);
			  DOPA_OUT : out  STD_LOGIC_VECTOR(3 downto 0);
			  ENB_IN : in STD_LOGIC;
           ADDRB_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DIB_IN : in  STD_LOGIC_VECTOR(31 downto 0);
			  DIPB_IN : in  STD_LOGIC_VECTOR(3 downto 0));
end BRAMHandler_CurveA_B00;

architecture Behavioral of BRAMHandler_CurveA_B00 is

	signal REGCEA: STD_LOGIC := '0';
	signal RSTA: STD_LOGIC := '0';
	signal WEA : STD_LOGIC_VECTOR(3 downto 0)  := (others => '0');
	signal DIA : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DIPA : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');

	signal DOB : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DOPB : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');
	signal REGCEB: STD_LOGIC := '0';
	signal RSTB: STD_LOGIC := '0';
	signal WEB : STD_LOGIC_VECTOR(3 downto 0) := (others => '1');
	
begin

	-- RAMB16BWER: 16k-bit Data and 2k-bit Parity Configurable Synchronous Dual Port Block RAM with Optional Output Registers
   --             Spartan-6
   -- Xilinx HDL Language Template, version 14.7

   RAMB16BWER_inst00 : RAMB16BWER
   generic map (
      -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
      DATA_WIDTH_A => DataWidth,
      DATA_WIDTH_B => DataWidth,
      -- DOA_REG/DOB_REG: Optional output register (0 or 1)
      DOA_REG => 0,
      DOB_REG => 0,
      -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
      EN_RSTRAM_A => TRUE,
      EN_RSTRAM_B => TRUE,
     	-- INITP_00 to INITP_07: Initial memory contents.
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

		-- INIT_00 to INIT_3F: Initial memory contents.
		INIT_00 => X"02F202BF028D025B022901F601C40192015F012D00FB00C90096006400320000",
		INIT_01 => X"061505E305B1057F054D051A04E804B604840451041F03ED03BB038803560324",
		INIT_02 => X"0938090608D408A20870083E080B07D907A707750743071106DE06AC067A0648",
		INIT_03 => X"0C5A0C280BF60BC40B920B600B2E0AFC0AC90A970A650A330A0109CF099D096B",
		INIT_04 => X"0F7A0F480F160EE40EB20E800E4E0E1C0DEA0DB80D860D540D220CF00CBE0C8C",
		INIT_05 => X"129712651233120211D0119E116C113A110910D710A510731041100F0FDD0FAC",
		INIT_06 => X"15B11580154E151D14EB14B914881456142413F313C1138F135E132C12FA12C9",
		INIT_07 => X"18C8189718661834180317D117A0176F173D170C16DA16A916771646161415E3",
		INIT_08 => X"1BDB1BAA1B791B481B171AE61AB51A841A521A2119F019BF198D195C192B18FA",
		INIT_09 => X"1EEA1EBA1E891E581E271DF61DC51D941D631D331D021CD11CA01C6F1C3E1C0D",
		INIT_0A => X"21F421C4219421632132210220D120A12070203F200F1FDE1FAD1F7D1F4C1F1B",
		INIT_0B => X"24F924C9249924692439240823D823A823782347231722E722B6228622552225",
		INIT_0C => X"27F927C9279927692739270926DA26AA267A264A261A25EA25BA258A255A252A",
		INIT_0D => X"2AF22AC22A932A632A342A0429D529A529762946291728E728B7288828582828",
		INIT_0E => X"2DE42DB52D862D572D282CF92CCA2C9B2C6C2C3D2C0D2BDE2BAF2B802B502B21",
		INIT_0F => X"30CF30A13072304430152FE72FB82F892F5B2F2C2EFD2ECE2EA02E712E422E13",
		INIT_10 => X"33B333853357332932FB32CD329F32703242321431E631B73189315B312C30FE",
		INIT_11 => X"368F36613634360635D935AB357D3550352234F434C73499346B343D340F33E1",
		INIT_12 => X"39623935390838DB38AE38813854382737FA37CC379F37723745371736EA36BC",
		INIT_13 => X"3C2D3C003BD43BA83B7B3B4F3B223AF53AC93A9C3A6F3A433A1639E939BC398F",
		INIT_14 => X"3EEE3EC23E963E6B3E3F3E133DE73DBB3D8F3D633D363D0A3CDE3CB23C863C59",
		INIT_15 => X"41A6417A414F412440F940CD40A24077404B40203FF43FC93F9D3F713F463F1A",
		INIT_16 => X"4453442943FE43D343A9437E4353432842FE42D342A8427D4252422741FC41D1",
		INIT_17 => X"46F646CC46A24678464E462445FA45D045A6457C4551452744FD44D244A8447E",
		INIT_18 => X"498E4965493C491248E948C04896486D4843481A47F047C7479D4773474A4720",
		INIT_19 => X"4C1A4BF24BCA4BA14B784B504B274AFE4AD64AAD4A844A5B4A324A0949E049B7",
		INIT_1A => X"4E9B4E744E4C4E244DFC4DD44DAC4D844D5C4D344D0C4CE44CBC4C944C6B4C43",
		INIT_1B => X"511050E950C2509B5074504D50264FFE4FD74FB04F894F614F3A4F124EEB4EC3",
		INIT_1C => X"53785352532C530652DF52B95293526C5246521F51F951D251AB5185515E5137",
		INIT_1D => X"55D455AE55895563553E551854F354CD54A85482545C5436541053EA53C4539E",
		INIT_1E => X"582257FD57D957B4578F576B5746572156FC56D756B2568D56685643561E55F9",
		INIT_1F => X"5A625A3F5A1B59F759D359AF598C59685944592058FB58D758B3588F586A5846",
		INIT_20 => X"5C955C725C4F5C2C5C095BE65BC35BA05B7D5B5A5B375B135AF05ACD5AA95A86",
		INIT_21 => X"5EB95E975E755E535E315E0F5DED5DCB5DA95D865D645D425D1F5CFD5CDA5CB7",
		INIT_22 => X"60CF60AE608D606C604B602960085FE75FC65FA45F835F615F405F1E5EFC5EDB",
		INIT_23 => X"62D562B56295627562556235621561F461D461B36193617261526131611060EF",
		INIT_24 => X"64CD64AE648F647064506431641263F263D363B36394637463556335631562F5",
		INIT_25 => X"66B566976679665A663C661E660065E165C365A46586656765486529650B64EC",
		INIT_26 => X"688D687068536835681867FB67DE67C067A367856768674A672C670E66F166D3",
		INIT_27 => X"6A556A396A1D6A0069E469C869AC698F69736956693A691D690068E368C768AA",
		INIT_28 => X"6C0C6BF16BD66BBB6BA06B856B696B4E6B336B176AFB6AE06AC46AA86A8D6A71",
		INIT_29 => X"6DB36D996D7F6D656D4B6D316D166CFC6CE26CC76CAD6C926C776C5D6C426C27",
		INIT_2A => X"6F496F306F176EFE6EE56ECC6EB36E9A6E806E676E4D6E346E1A6E006DE76DCD",
		INIT_2B => X"70CE70B6709E7086706E7056703E7026700E6FF56FDD6FC46FAC6F936F7B6F62",
		INIT_2C => X"7241722A721471FD71E671CF71B871A1718A7172715B7144712C711570FD70E5",
		INIT_2D => X"73A3738D73787362734C73367320730A72F472DE72C872B2729B7285726E7258",
		INIT_2E => X"74F374DE74CA74B574A0748C74777462744D74387423740E73F973E373CE73B8",
		INIT_2F => X"7631761D760A75F675E375CF75BC75A875947580756C755875447530751B7507",
		INIT_30 => X"775C774A773877257713770176EE76DB76C976B676A37690767D766A76577644",
		INIT_31 => X"787578647853784278317820780E77FD77EB77DA77C877B677A477927780776E",
		INIT_32 => X"797C796C795C794C793C792C791C790B78FB78EB78DA78C978B978A878977886",
		INIT_33 => X"7A707A617A527A447A357A267A177A0879F879E979DA79CA79BB79AB799C798C",
		INIT_34 => X"7B517B437B367B287B1A7B0D7AFF7AF17AE37AD57AC77AB87AAA7A9C7A8D7A7F",
		INIT_35 => X"7C1F7C137C067BFA7BED7BE17BD47BC77BBA7BAD7BA07B937B867B797B6C7B5E",
		INIT_36 => X"7CDA7CCF7CC37CB87CAD7CA17C967C8A7C7F7C737C677C5B7C4F7C437C377C2B",
		INIT_37 => X"7D817D777D6D7D637D597D4F7D457D3A7D307D257D1B7D107D057CFB7CF07CE5",
		INIT_38 => X"7E157E0D7E047DFB7DF27DE97DE07DD77DCE7DC47DBB7DB27DA87D9E7D957D8B",
		INIT_39 => X"7E967E8F7E877E7F7E787E707E687E607E587E507E487E407E377E2F7E277E1E",
		INIT_3A => X"7F037EFD7EF77EF07EEA7EE37EDD7ED67ECF7EC87EC17EBA7EB37EAC7EA57E9E",
		INIT_3B => X"7F5D7F587F537F4E7F487F437F3E7F387F337F2D7F277F217F1C7F167F107F09",
		INIT_3C => X"7FA37F9F7F9B7F977F937F8F7F8B7F877F827F7E7F797F757F707F6C7F677F62",
		INIT_3D => X"7FD57FD37FD07FCD7FCA7FC87FC57FC27FBE7FBB7FB87FB57FB17FAE7FAA7FA7",
		INIT_3E => X"7FF47FF27FF17FEF7FEE7FEC7FEB7FE97FE77FE57FE37FE17FDF7FDC7FDA7FD8",
		INIT_3F => X"7FFE7FFE7FFE7FFE7FFE7FFD7FFD7FFC7FFC7FFB7FFA7FF97FF87FF77FF67FF5",
      -- INIT_A/INIT_B: Initial values on output port
      INIT_A => X"000000000",
      INIT_B => X"000000000",
      -- INIT_FILE: Optional file used to specify initial RAM contents
      INIT_FILE => "NONE",
      -- RSTTYPE: "SYNC" or "ASYNC" 
      RSTTYPE => "SYNC",
      -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
      RST_PRIORITY_A => "CE",
      RST_PRIORITY_B => "CE",
      -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
      SIM_COLLISION_CHECK => "ALL",
      -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
      SIM_DEVICE => "SPARTAN6",
      -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
      SRVAL_A => X"000000000",
      SRVAL_B => X"000000000",
      -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
      WRITE_MODE_A => "READ_FIRST",
      WRITE_MODE_B => "READ_FIRST" 
   )
   port map (
      -- Port A Data: 32-bit (each) output: Port A data
      DOA => DOA_OUT,       -- 32-bit output: A port data output
      DOPA => DOPA_OUT,     -- 4-bit output: A port parity output
      -- Port B Data: 32-bit (each) output: Port B data
      DOB => DOB,       -- 32-bit output: B port data output
      DOPB => DOPB,     -- 4-bit output: B port parity output
      -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
      ADDRA => ADDRA_IN,   -- 14-bit input: A port address input
      CLKA => CLK_IN,     -- 1-bit input: A port clock input
      ENA => ENA_IN,       -- 1-bit input: A port enable input
      REGCEA => REGCEA, -- 1-bit input: A port register clock enable input
      RSTA => RSTA,     -- 1-bit input: A port register set/reset input
      WEA => WEA,       -- 4-bit input: Port A byte-wide write enable input
      -- Port A Data: 32-bit (each) input: Port A data
      DIA => DIA,       -- 32-bit input: A port data input
      DIPA => DIPA,     -- 4-bit input: A port parity input
      -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
      ADDRB => ADDRB_IN,   -- 14-bit input: B port address input
      CLKB => CLK_IN,     -- 1-bit input: B port clock input
      ENB => ENB_IN,       -- 1-bit input: B port enable input
      REGCEB => REGCEB, -- 1-bit input: B port register clock enable input
      RSTB => RSTB,     -- 1-bit input: B port register set/reset input
      WEB => WEB,       -- 4-bit input: Port B byte-wide write enable input
      -- Port B Data: 32-bit (each) input: Port B data
      DIB => DIB_IN,       -- 32-bit input: B port data input
      DIPB => DIPB_IN      -- 4-bit input: B port parity input
   );
	
   -- End of RAMB16BWER_inst instantiation
end Behavioral;

