----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:07:53 11/05/2021 
-- Design Name: 
-- Module Name:    BRAMHandler - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity BRAMHandler_CurveB_B11 is
	 Generic ( DataWidth : integer := 18);
    Port ( CLK_IN : in  STD_LOGIC;
			  ENA_IN : in STD_LOGIC;
           ADDRA_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DOA_OUT : out  STD_LOGIC_VECTOR(31 downto 0);
			  DOPA_OUT : out  STD_LOGIC_VECTOR(3 downto 0);
			  ENB_IN : in STD_LOGIC;
           ADDRB_IN : in  STD_LOGIC_VECTOR(13 downto 0);
           DIB_IN : in  STD_LOGIC_VECTOR(31 downto 0);
			  DIPB_IN : in  STD_LOGIC_VECTOR(3 downto 0));
end BRAMHandler_CurveB_B11;

architecture Behavioral of BRAMHandler_CurveB_B11 is

	signal REGCEA: STD_LOGIC := '0';
	signal RSTA: STD_LOGIC := '0';
	signal WEA : STD_LOGIC_VECTOR(3 downto 0)  := (others => '0');
	signal DIA : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DIPA : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');

	signal DOB : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
	signal DOPB : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');
	signal REGCEB: STD_LOGIC := '0';
	signal RSTB: STD_LOGIC := '0';
	signal WEB : STD_LOGIC_VECTOR(3 downto 0) := (others => '1');
	
begin

	-- RAMB16BWER: 16k-bit Data and 2k-bit Parity Configurable Synchronous Dual Port Block RAM with Optional Output Registers
   --             Spartan-6
   -- Xilinx HDL Language Template, version 14.7

   RAMB16BWER_inst11 : RAMB16BWER
   generic map (
      -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
      DATA_WIDTH_A => DataWidth,
      DATA_WIDTH_B => DataWidth,
      -- DOA_REG/DOB_REG: Optional output register (0 or 1)
      DOA_REG => 0,
      DOB_REG => 0,
      -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
      EN_RSTRAM_A => TRUE,
      EN_RSTRAM_B => TRUE,
      -- INITP_00 to INITP_07: Initial memory contents.
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

		-- INIT_00 to INIT_3F: Initial memory contents.
		INIT_00 => X"C006C006C005C005C004C004C003C003C003C002C002C002C002C002C002C002",
		INIT_01 => X"C015C014C013C011C010C00FC00EC00DC00CC00BC00BC00AC009C008C008C007",
		INIT_02 => X"C02DC02CC02AC028C026C025C023C022C020C01EC01DC01CC01AC019C017C016",
		INIT_03 => X"C050C04DC04BC049C046C044C042C040C03DC03BC039C037C035C033C031C02F",
		INIT_04 => X"C07CC079C076C073C070C06DC06AC067C065C062C05FC05DC05AC057C055C052",
		INIT_05 => X"C0B2C0AEC0ABC0A7C0A4C0A0C09DC099C096C092C08FC08CC089C085C082C07F",
		INIT_06 => X"C0F2C0EDC0E9C0E5C0E1C0DDC0D9C0D5C0D1C0CDC0C9C0C5C0C1C0BDC0B9C0B6",
		INIT_07 => X"C13BC136C132C12DC128C123C11FC11AC115C111C10CC108C103C0FFC0FAC0F6",
		INIT_08 => X"C18EC189C183C17EC179C173C16EC169C164C15EC159C154C14FC14AC145C140",
		INIT_09 => X"C1EBC1E5C1DFC1D9C1D3C1CDC1C7C1C1C1BCC1B6C1B0C1AAC1A5C19FC199C194",
		INIT_0A => X"C252C24BC244C23EC237C231C22AC224C21DC217C210C20AC204C1FEC1F7C1F1",
		INIT_0B => X"C2C1C2BAC2B3C2ACC2A5C29DC296C28FC288C281C27AC274C26DC266C25FC258",
		INIT_0C => X"C33BC333C32BC323C31CC314C30CC305C2FDC2F5C2EEC2E6C2DFC2D7C2D0C2C9",
		INIT_0D => X"C3BEC3B5C3ADC3A4C39CC394C38BC383C37BC373C36BC363C35BC353C34BC343",
		INIT_0E => X"C44AC441C438C42FC426C41DC414C40BC402C3FAC3F1C3E8C3E0C3D7C3CFC3C6",
		INIT_0F => X"C4DFC4D5C4CCC4C2C4B9C4AFC4A6C49CC493C48AC480C477C46EC465C45CC453",
		INIT_10 => X"C57DC573C569C55FC555C54BC541C537C52DC523C519C50FC506C4FCC4F2C4E8",
		INIT_11 => X"C625C61AC60FC604C5FAC5EFC5E5C5DAC5D0C5C5C5BBC5B0C5A6C59CC592C587",
		INIT_12 => X"C6D5C6CAC6BEC6B3C6A8C69DC692C687C67CC671C666C65BC650C645C63AC62F",
		INIT_13 => X"C78EC782C776C76BC75FC753C747C73CC730C725C719C70EC702C6F7C6EBC6E0",
		INIT_14 => X"C850C843C837C82BC81FC812C806C7FAC7EEC7E2C7D6C7CAC7BEC7B2C7A6C79A",
		INIT_15 => X"C91AC90DC900C8F4C8E7C8DAC8CDC8C1C8B4C8A7C89BC88EC882C875C869C85C",
		INIT_16 => X"C9EDC9E0C9D2C9C5C9B8C9AAC99DC990C983C975C968C95BC94EC941C934C927",
		INIT_17 => X"CAC8CABACAACCA9FCA91CA83CA75CA67CA5ACA4CCA3ECA31CA23CA16CA08C9FB",
		INIT_18 => X"CBACCB9DCB8FCB81CB72CB64CB56CB47CB39CB2BCB1DCB0FCB00CAF2CAE4CAD6",
		INIT_19 => X"CC97CC88CC79CC6BCC5CCC4DCC3ECC2FCC21CC12CC03CBF5CBE6CBD7CBC9CBBA",
		INIT_1A => X"CD8BCD7BCD6CCD5DCD4DCD3ECD2FCD1FCD10CD01CCF2CCE3CCD3CCC4CCB5CCA6",
		INIT_1B => X"CE86CE76CE66CE56CE46CE37CE27CE17CE07CDF8CDE8CDD8CDC9CDB9CDAACD9A",
		INIT_1C => X"CF89CF79CF68CF58CF47CF37CF27CF17CF07CEF6CEE6CED6CEC6CEB6CEA6CE96",
		INIT_1D => X"D093D082D072D061D050D03FD02FD01ED00DCFFDCFECCFDBCFCBCFBACFAACF99",
		INIT_1E => X"D1A5D194D182D171D160D14FD13DD12CD11BD10AD0F9D0E8D0D7D0C6D0B5D0A4",
		INIT_1F => X"D2BED2ACD29AD289D277D265D254D242D230D21FD20DD1FCD1EAD1D9D1C8D1B6",
		INIT_20 => X"D3DED3CBD3B9D3A7D395D383D371D35FD34DD33BD329D317D305D2F3D2E1D2D0",
		INIT_21 => X"D504D4F2D4DFD4CCD4BAD4A7D495D482D470D45ED44BD439D427D414D402D3F0",
		INIT_22 => X"D631D61ED60BD5F8D5E5D5D3D5C0D5ADD59AD587D574D562D54FD53CD529D517",
		INIT_23 => X"D765D752D73ED72BD718D704D6F1D6DED6CAD6B7D6A4D691D67ED66BD658D644",
		INIT_24 => X"D89FD88BD877D864D850D83CD829D815D801D7EED7DAD7C7D7B3D7A0D78CD779",
		INIT_25 => X"D9DFD9CBD9B7D9A3D98FD97AD966D952D93ED92AD916D902D8EFD8DBD8C7D8B3",
		INIT_26 => X"DB25DB10DAFCDAE7DAD3DABFDAAADA96DA81DA6DDA59DA44DA30DA1CDA08D9F3",
		INIT_27 => X"DC71DC5CDC47DC32DC1DDC08DBF4DBDFDBCADBB5DBA1DB8CDB77DB63DB4EDB3A",
		INIT_28 => X"DDC2DDADDD97DD82DD6DDD58DD43DD2EDD19DD03DCEEDCD9DCC4DCAFDC9ADC86",
		INIT_29 => X"DF18DF03DEEDDED8DEC2DEADDE97DE82DE6CDE57DE42DE2CDE17DE02DDECDDD7",
		INIT_2A => X"E074E05EE048E032E01CE006DFF1DFDBDFC5DFB0DF9ADF84DF6EDF59DF43DF2E",
		INIT_2B => X"E1D4E1BEE1A8E191E17BE165E14FE139E123E10DE0F7E0E1E0CBE0B5E09FE089",
		INIT_2C => X"E339E322E30CE2F6E2DFE2C9E2B2E29CE286E26FE259E243E22DE216E200E1EA",
		INIT_2D => X"E4A2E48CE475E45EE448E431E41AE404E3EDE3D6E3C0E3A9E393E37CE366E34F",
		INIT_2E => X"E610E5F9E5E2E5CBE5B4E59DE586E56FE559E542E52BE514E4FDE4E7E4D0E4B9",
		INIT_2F => X"E782E76AE753E73CE725E70EE6F6E6DFE6C8E6B1E69AE683E66CE655E63EE627",
		INIT_30 => X"E8F7E8E0E8C8E8B1E899E882E86BE853E83CE824E80DE7F6E7DFE7C7E7B0E799",
		INIT_31 => X"EA70EA58EA41EA29EA11E9FAE9E2E9CBE9B3E99BE984E96CE955E93DE926E90E",
		INIT_32 => X"EBECEBD4EBBDEBA5EB8DEB75EB5DEB45EB2EEB16EAFEEAE6EACFEAB7EA9FEA88",
		INIT_33 => X"ED6CED54ED3CED24ED0CECF4ECDCECC4ECACEC94EC7CEC64EC4CEC34EC1CEC04",
		INIT_34 => X"EEEEEED6EEBDEEA5EE8DEE75EE5DEE45EE2CEE14EDFCEDE4EDCCEDB4ED9CED84",
		INIT_35 => X"F073F05AF042F02AF011EFF9EFE1EFC8EFB0EF98EF7FEF67EF4FEF37EF1EEF06",
		INIT_36 => X"F1FAF1E2F1C9F1B1F198F180F167F14FF136F11EF105F0EDF0D4F0BCF0A4F08B",
		INIT_37 => X"F384F36BF352F33AF321F308F2F0F2D7F2BFF2A6F28DF275F25CF244F22BF213",
		INIT_38 => X"F50FF4F6F4DDF4C5F4ACF493F47AF462F449F430F418F3FFF3E6F3CEF3B5F39C",
		INIT_39 => X"F69CF683F66AF651F639F620F607F5EEF5D5F5BCF5A4F58BF572F559F541F528",
		INIT_3A => X"F82BF812F7F9F7E0F7C7F7AEF795F77CF763F74AF731F718F700F6E7F6CEF6B5",
		INIT_3B => X"F9BAF9A1F988F96FF956F93DF924F90BF8F2F8D9F8C0F8A7F88EF875F85CF844",
		INIT_3C => X"FB4BFB32FB19FB00FAE7FACEFAB5FA9CFA83FA69FA50FA37FA1EFA05F9ECF9D3",
		INIT_3D => X"FCDCFCC3FCAAFC91FC78FC5FFC46FC2DFC14FBFBFBE1FBC8FBAFFB96FB7DFB64",
		INIT_3E => X"FE6EFE55FE3CFE23FE0AFDF1FDD8FDBEFDA5FD8CFD73FD5AFD41FD28FD0FFCF6",
		INIT_3F => X"0000FFE7FFCEFFB5FF9CFF83FF6AFF51FF37FF1EFF05FEECFED3FEBAFEA1FE87",
      -- INIT_A/INIT_B: Initial values on output port
      INIT_A => X"000000000",
      INIT_B => X"000000000",
      -- INIT_FILE: Optional file used to specify initial RAM contents
      INIT_FILE => "NONE",
      -- RSTTYPE: "SYNC" or "ASYNC" 
      RSTTYPE => "SYNC",
      -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
      RST_PRIORITY_A => "CE",
      RST_PRIORITY_B => "CE",
      -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
      SIM_COLLISION_CHECK => "ALL",
      -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
      SIM_DEVICE => "SPARTAN6",
      -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
      SRVAL_A => X"000000000",
      SRVAL_B => X"000000000",
      -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
      WRITE_MODE_A => "READ_FIRST",
      WRITE_MODE_B => "READ_FIRST" 
   )
   port map (
      -- Port A Data: 32-bit (each) output: Port A data
      DOA => DOA_OUT,       -- 32-bit output: A port data output
      DOPA => DOPA_OUT,     -- 4-bit output: A port parity output
      -- Port B Data: 32-bit (each) output: Port B data
      DOB => DOB,       -- 32-bit output: B port data output
      DOPB => DOPB,     -- 4-bit output: B port parity output
      -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
      ADDRA => ADDRA_IN,   -- 14-bit input: A port address input
      CLKA => CLK_IN,     -- 1-bit input: A port clock input
      ENA => ENA_IN,       -- 1-bit input: A port enable input
      REGCEA => REGCEA, -- 1-bit input: A port register clock enable input
      RSTA => RSTA,     -- 1-bit input: A port register set/reset input
      WEA => WEA,       -- 4-bit input: Port A byte-wide write enable input
      -- Port A Data: 32-bit (each) input: Port A data
      DIA => DIA,       -- 32-bit input: A port data input
      DIPA => DIPA,     -- 4-bit input: A port parity input
      -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
      ADDRB => ADDRB_IN,   -- 14-bit input: B port address input
      CLKB => CLK_IN,     -- 1-bit input: B port clock input
      ENB => ENB_IN,       -- 1-bit input: B port enable input
      REGCEB => REGCEB, -- 1-bit input: B port register clock enable input
      RSTB => RSTB,     -- 1-bit input: B port register set/reset input
      WEB => WEB,       -- 4-bit input: Port B byte-wide write enable input
      -- Port B Data: 32-bit (each) input: Port B data
      DIB => DIB_IN,       -- 32-bit input: B port data input
      DIPB => DIPB_IN      -- 4-bit input: B port parity input
   );


   -- End of RAMB16BWER_inst instantiation
end Behavioral;

